-- -------------------------------------------------------
-- The files contains UART Transmitter architecture.
-- Author :- Rishi Vaghasiya (35869)
-- Wintersemester 2023/24
-- -------------------------------------------------------

architecture of rv_UART_TX_a of rv_UART_TX_e is 
end rv_UART_TX_a;
